module ex;
assign y=a&b;
endmodule

